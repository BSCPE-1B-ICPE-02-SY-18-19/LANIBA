CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 4 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
110100498 0
0
6 Title:
5 Name:
0
0
0
12
5 SAVE-
218 414 378 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
5130 0 0
2
5.89884e-315 0
0
7 Ground~
168 1144 271 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
391 0 0
2
5.89884e-315 5.26354e-315
0
6 74112~
219 938 314 0 7 32
0 6 4 3 4 6 18 17
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U1B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 5 0
1 U
3124 0 0
2
5.89884e-315 5.30499e-315
0
6 74112~
219 736 315 0 7 32
0 6 5 3 5 6 19 16
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 5 0
1 U
3421 0 0
2
5.89884e-315 5.32571e-315
0
6 74112~
219 523 315 0 7 32
0 6 7 3 7 6 20 15
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U5B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 4 0
1 U
8157 0 0
2
5.89884e-315 5.34643e-315
0
6 74112~
219 307 315 0 7 32
0 6 6 3 6 6 21 7
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U5A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 4 0
1 U
5572 0 0
2
5.89884e-315 5.3568e-315
0
9 2-In AND~
219 829 222 0 3 22
0 5 16 4
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
8901 0 0
2
5.89884e-315 5.36716e-315
0
9 2-In AND~
219 629 214 0 3 22
0 7 15 5
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7361 0 0
2
5.89884e-315 5.37752e-315
0
2 +V
167 307 199 0 1 3
0 6
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4747 0 0
2
5.89884e-315 5.38788e-315
0
9 CC 7-Seg~
183 1060 309 0 17 19
10 14 13 12 11 10 9 8 22 2
0 0 1 1 1 1 1 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
972 0 0
2
5.89884e-315 5.39306e-315
0
6 74LS48
188 1023 489 0 14 29
0 17 16 15 7 23 24 8 9 10
11 12 13 14 25
0
0 0 4832 0
7 74LS248
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3472 0 0
2
5.89884e-315 5.39824e-315
0
7 Pulser~
4 160 290 0 10 12
0 26 27 28 3 0 0 5 5 4
8
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9998 0 0
2
5.89884e-315 5.40342e-315
0
36
4 0 0 0 0 0 0 12 0 0 14 5
190 290
190 324
246 324
246 378
251 378
9 1 2 0 0 8320 0 10 2 0 0 4
1060 267
1060 163
1144 163
1144 265
0 3 3 0 0 4096 0 0 3 13 0 4
703 378
899 378
899 287
908 287
4 2 4 0 0 4096 0 3 3 0 0 4
914 296
891 296
891 278
914 278
0 0 5 0 0 4096 0 0 0 21 6 3
684 279
650 279
650 180
3 1 5 0 0 4224 0 8 7 0 0 5
650 214
650 180
650 180
650 213
805 213
0 0 6 0 0 4096 0 0 0 8 19 2
405 244
405 332
0 0 6 0 0 4096 0 0 0 9 16 2
307 244
523 244
0 0 6 0 0 0 0 0 0 23 10 3
260 279
260 244
307 244
1 1 6 0 0 0 0 9 6 0 0 2
307 208
307 252
0 1 7 0 0 12288 0 0 8 12 0 4
476 279
443 279
443 205
605 205
4 0 7 0 0 0 0 5 0 0 31 3
499 297
476 297
476 279
0 3 3 0 0 0 0 0 4 14 0 4
485 378
703 378
703 288
706 288
3 3 3 0 0 12416 0 6 5 0 0 6
277 288
251 288
251 378
485 378
485 288
493 288
0 1 6 0 0 0 0 0 3 16 0 3
737 244
938 244
938 251
1 1 6 0 0 0 0 5 4 0 0 6
523 252
523 244
737 244
737 244
736 244
736 252
0 5 6 0 0 0 0 0 3 18 0 3
737 332
938 332
938 326
0 5 6 0 0 0 0 0 4 19 0 5
524 332
737 332
737 332
736 332
736 327
5 5 6 0 0 8320 0 6 5 0 0 6
307 327
307 332
524 332
524 332
523 332
523 327
0 3 4 0 0 8320 0 0 7 4 0 4
891 279
847 279
847 222
850 222
4 2 5 0 0 0 0 4 4 0 0 4
712 297
684 297
684 279
712 279
7 0 7 0 0 0 0 6 0 0 31 2
331 279
369 279
4 2 6 0 0 0 0 6 6 0 0 6
283 297
260 297
260 277
258 277
258 279
283 279
7 7 8 0 0 4224 0 10 11 0 0 5
1075 345
1075 397
1147 397
1147 453
1055 453
6 8 9 0 0 4224 0 10 11 0 0 5
1069 345
1069 402
1142 402
1142 462
1055 462
5 9 10 0 0 4224 0 10 11 0 0 5
1063 345
1063 407
1137 407
1137 471
1055 471
4 10 11 0 0 4224 0 10 11 0 0 5
1057 345
1057 412
1132 412
1132 480
1055 480
3 11 12 0 0 4224 0 10 11 0 0 5
1051 345
1051 417
1127 417
1127 489
1055 489
2 12 13 0 0 4224 0 10 11 0 0 5
1045 345
1045 422
1122 422
1122 498
1055 498
1 13 14 0 0 4224 0 10 11 0 0 5
1039 345
1039 427
1117 427
1117 507
1055 507
2 4 7 0 0 12416 0 5 11 0 0 4
499 279
369 279
369 480
991 480
0 3 15 0 0 8320 0 0 11 36 0 3
585 276
585 471
991 471
0 2 16 0 0 8320 0 0 11 35 0 3
793 276
793 462
991 462
7 1 17 0 0 8320 0 3 11 0 0 4
962 278
990 278
990 453
991 453
7 2 16 0 0 0 0 4 7 0 0 4
760 279
793 279
793 231
805 231
7 2 15 0 0 0 0 5 8 0 0 4
547 279
585 279
585 223
605 223
7
-27 0 0 0 400 0 0 0 0 3 2 1 34
14 Britannic Bold
0 0 0 14
928 21 1161 63
940 29 1148 59
14 MARCH 06, 2019
-37 0 0 0 700 0 0 0 0 3 2 1 82
8 Broadway
0 0 0 32
172 89 997 147
186 97 982 139
32 BINARY 4-BIT SYNCHRONOUS COUNTER
-19 0 0 0 400 0 0 0 0 3 2 1 34
14 Britannic Bold
0 0 0 8
32 42 138 71
43 50 126 71
8 BSCPE-1B
-24 0 0 0 700 0 0 0 0 3 2 1 18
20 Bernard MT Condensed
0 0 0 22
630 529 911 567
643 537 897 565
22 ENGR. MAX ANGELO PERIN
-16 0 0 0 400 255 0 0 0 3 2 1 66
15 Brush Script MT
0 0 0 13
489 510 626 539
500 518 614 537
13 SUBMITTED TO:
-16 0 0 0 400 255 0 0 0 3 2 1 66
15 Brush Script MT
0 0 0 13
9 512 146 541
20 520 134 539
13 SUBMITTED BY:
-27 0 0 0 400 0 0 0 0 3 2 1 34
14 Britannic Bold
0 0 0 21
141 522 453 564
153 530 440 560
21 LANIBA, ROTCHE MAE C.
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
